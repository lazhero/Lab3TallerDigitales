module Calc_test();

	logic [3:0] A,B,sel, Output;
	logic Z,O,Ca,Neg;
	ALU #(.N(4)) myALU (.A(A),.B(B),.sel(sel), .out(Output), .Z(Z),.O(O),.Ca(Ca),.Neg(Neg));
	initial begin 
	sel=4'b0000;
	A=4'b0011;
	B=4'b1101;
	#1;
	assert(Output==4'b1010) else $error("La suma falla");
	assert(Neg == 1)else $error("Bandera Neg falla sum");
	assert(Ca == 0)else $error("Bandera Carry falla sum");
	assert(Z == 0)else $error("Bandera Zero falla sum");
	assert(O == 0)else $error("Bandera Over falla sum");
	#1;

	sel=4'b0001;
	A=4'b0010;
	B=4'b1101;
	#1;
	assert(Output==4'b0111) else $error("La resta falla");
   assert(Neg == 0)else $error("Bandera Neg falla res");
	assert(Ca == 1)else $error("Bandera Carry falla res");
	assert(Z == 0)else $error("Bandera Zero falla res");
	assert(O == 0)else $error("Bandera Over falla res");
	#1;
	
	sel=4'b0010;
	A=4'b0011;
	B=4'b1001;
   #1;
	assert(Output==4'b1011) else $error("La multiplicacion falla");
	assert(Neg == 1)else $error("Bandera Neg falla mult");
	assert(Ca == 0)else $error("Bandera Carry falla mult");
	assert(Z == 0)else $error("Bandera Zero falla mult");
	assert(O == 1)else $error("Bandera Over falla mult");
	#1;
	sel=4'b0011;
	A=4'b0110;
	B=4'b1011;
	#1;
	assert(Output==4'b1010) else $error("La div falla");
	assert(Neg == 1)else $error("Bandera Neg falla div");
	assert(Ca == 0)else $error("Bandera Carry falla div");
	assert(Z == 0)else $error("Bandera Zero falla div");
	assert(O == 0)else $error("Bandera Over falla div");
	#1;
	sel=4'b0100;
	A=4'b0011;
	B=4'b0001;
	#1;
	assert(Output==4'b0000) else $error("el mod falla");
	assert(Neg == 0)else $error("Bandera Neg falla mod");
	assert(Ca == 0)else $error("Bandera Carry falla mod");
	assert(Z == 1)else $error("Bandera Zero falla mod");
	assert(O == 0)else $error("Bandera Over falla mod");
	#1;
	sel=4'b0101;
	A=4'b0010;
	B=4'b0001;
	#1;
	assert(Output==4'b0100) else $error("La ShiftL falla");
   assert(Neg == 0)else $error("Bandera Neg falla ShiftL");
	assert(Ca == 0)else $error("Bandera Carry falla ShiftL");
	assert(Z == 0)else $error("Bandera Zero falla ShiftL");
	assert(O == 0)else $error("Bandera Over falla ShiftL");
	#1;
	sel=4'b0110;
	A=4'b0011;
	B=4'b0001;
	#1;
	assert(Output==4'b0001) else $error("La ShiftR falla");
	assert(Neg == 0)else $error("Bandera Neg falla ShiftR");
	assert(Ca == 0)else $error("Bandera Carry falla ShiftR");
	assert(Z == 0)else $error("Bandera Zero falla ShiftR");
	assert(O == 0)else $error("Bandera Over falla ShiftR");
	#1;
	sel=4'b0111;
	A=4'b0110;
	B=4'b1011;
	#1;
	assert(Output==4'b0010) else $error("La And falla");
	assert(Neg == 0)else $error("Bandera Neg falla And");
	assert(Ca == 0)else $error("Bandera Carry falla And");
	assert(Z == 0)else $error("Bandera Zero falla And");
	assert(O == 0)else $error("Bandera Over falla And");
	#1;
	sel=4'b1001;
	A=4'b0110;
	B=4'b1011;
	
	#1;
	assert(Output==4'b1111) else $error("La OR falla");
	assert(Neg == 1)else $error("Bandera Neg falla OR");
	assert(Ca == 0)else $error("Bandera Carry falla OR");
	assert(Z == 0)else $error("Bandera Zero falla OR");
	assert(O == 0)else $error("Bandera Over falla OR");
	#1;
	sel=4'b1000;
	A=4'b0110;
	B=4'b1011;
	#1;
	assert(Output==4'b1101) else $error("La XOR falla");
	assert(Neg == 1)else $error("Bandera Neg falla XOR");
	assert(Ca == 0)else $error("Bandera Carry falla XOR");
	assert(Z == 0)else $error("Bandera Zero falla XOR");
	assert(O == 0)else $error("Bandera Over falla XOR");
	#1;
	end
endmodule 